altfp_convert_int_to_float_inst : altfp_convert_int_to_float PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
