altfp_convert_float_to_int_inst : altfp_convert_float_to_int PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
